`timescale 1ns / 1ps
/*******************************************************************
*
* Module: module_Instruction_Memory.v
* Project: Archetchture_project
* Author: Mariam Abulela     900141674
          Nada Badawy        900171975
          Mohamed Al-Awadly  900163100
* Description: in this module we get the address of the instruction
* that should be fetched in the instruction memory to have the instruction
* Change history: 03/10/19 � creat the module
* 28/10/19 � Edit the module 
*
**********************************************************************/

module Instmem (
input [11:0] address,
output [31:0] instruction);

 reg [7:0] mem [(4*1024-1):0];
 initial begin
 $readmemh("E:/Fall 19/arch/New folder/Branch.hex", mem); 
 end 
// initial begin
 
 
 
 
 
// mem[0]=8'b00000000;
// mem[1]=8'b0000_0000;
// mem[2]=8'b0_010_0000;
// mem[3]=8'b1_0000011; //lw x1, 0(x0)
// mem[4]=8'b0000000_0;
// mem[5]=8'b0000_0000;
// mem[6]=8'b0_000_0000;
// mem[7]=8'b0_0110011 ; //add x0, x0, x0
// mem[8]=8'b0000000_0;
// mem[9]=8'b0000_0000;
// mem[10]=8'b0_000_0000;
// mem[11]=8'b0_0110011 ; //add x0, x0, x0
// mem[12]=8'b0000000_0;
// mem[13]=8'b0000_0000;
 
// mem[14]=8'b0_000_0000;
// mem[15]=8'b0_0110011 ; //add x0, x0, x0
// mem[16]=8'b00000000;
// mem[17]=8'b0100_0000;
// mem[18]=8'b0_010_0001;
// mem[19]=8'b0_0000011 ; //lw x2, 4(x0)
// mem[20]=8'b0000000_0;
// mem[21]=8'b0000_0000;
// mem[22]=8'b0_000_0000;
// mem[23]=8'b0_0110011 ; //add x0, x0, x0
// mem[24]=8'b0000000_0;
// mem[25]=8'b0000_0000;
// mem[26]=8'b0_000_0000;
// mem[27]=8'b0_0110011 ; //add x0, x0, x0
// mem[28]=8'b0000000_0;
// mem[29]=8'b0000_0000;
// mem[30]=8'b0_000_0000;
// mem[31]=8'b0_0110011 ; //add x0, x0, x0
// mem[32]=8'b00000000;
// mem[33]=8'b1000_0000;
// mem[34]=8'b0_010_0001;
// mem[35]=8'b1_0000011 ; //lw x3, 8(x0)
// mem[36]=8'b0000000_0;
// mem[37]=8'b0000_0000;
// mem[38]=8'b0_000_0000;
// mem[39]=8'b0_0110011 ; //add x0, x0, x0
// mem[40]=8'b0000000_0;
// mem[41]=8'b0000_0000;
// mem[42]=8'b0_000_0000;
// mem[43]=8'b0_0110011 ; //add x0, x0, x0
// mem[44]=8'b0000000_0;
// mem[45]=8'b0000_0000;
// mem[46]=8'b0_000_0000;
// mem[47]=8'b0_0110011 ; //add x0, x0, x0
// mem[48]=8'b0000000_0;
// mem[49]=8'b0010_0000;
// mem[50]=8'b1_110_0010;
// mem[51]=8'b0_0110011 ; //or x4, x1, x2
// mem[52]=8'b0000000_0;
// mem[53]=8'b0000_0000;
// mem[54]=8'b0_000_0000;
// mem[55]=8'b0_0110011 ; //add x0, x0, x0
// mem[56]=8'b0000000_0;
// mem[57]=8'b0000_0000;
// mem[58]=8'b0_000_0000;
// mem[59]=8'b0_0110011 ; //add x0, x0, x0
// mem[60]=8'b0000000_0;
// mem[61]=8'b0000_0000;
// mem[62]=8'b0_000_0000;
// mem[63]=8'b0_0110011 ; //add x0, x0, x0
// mem[64]=8'b0_000001_0;
// mem[65]=8'b0011_0010;
// mem[66]=8'b0_000_0000;
// mem[67]=8'b_0_1100011; //beq x4, x3, 16
// mem[68]=8'b0000000_0;
// mem[69]=8'b0000_0000;
// mem[70]=8'b0_000_0000;
// mem[71]=8'b0_0110011 ; //add x0, x0, x0
// mem[72]=8'b0000000_0;
// mem[73]=8'b0000_0000;
// mem[74]=8'b0_000_0000;
// mem[75]=8'b0_0110011 ; //add x0, x0, x0
// mem[76]=8'b0000000_0;
// mem[77]=8'b0000_0000;
// mem[78]=8'b0_000_0000;
// mem[79]=8'b0_0110011 ; //add x0, x0, x0
// mem[80]=8'b0000000_0;
// mem[81]=8'b0010_0000;
// mem[82]=8'b1_000_0001;
// mem[83]=8'b1_0110011 ; //add x3, x1, x2
// mem[84]=8'b0000000_0;
// mem[85]=8'b0000_0000;
// mem[86]=8'b0_000_0000;
// mem[87]=8'b0_0110011 ; //add x0, x0, x0
// mem[88]=8'b0000000_0;
// mem[89]=8'b0000_0000;
// mem[90]=8'b0_000_0000;
// mem[91]=8'b0_0110011 ; //add x0, x0, x0
// mem[92]=8'b0000000_0;
// mem[93]=8'b0000_0000;
// mem[94]=8'b0_000_0000;
// mem[95]=8'b0_0110011 ; //add x0, x0, x0
// mem[96]=8'b0000000_0;
// mem[97]=8'b0010_0001;
// mem[98]=8'b1_000_0010;
// mem[99]=8'b1_0110011 ; //add x5, x3, x2
// mem[100]=8'b0000000_0;
// mem[101]=8'b0000_0000;
// mem[102]=8'b0_000_0000;
// mem[103]=8'b0_0110011 ; //add x0, x0, x0
// mem[104]=8'b0000000_0;
// mem[105]=8'b0000_0000;
// mem[106]=8'b0_000_0000;
// mem[107]=8'b0_0110011 ; //add x0, x0, x0
// mem[108]=8'b0000000_0;
// mem[109]=8'b0000_0000;
// mem[110]=8'b0_000_0000;
// mem[111]=8'b0_0110011 ; //add x0, x0, x0
// mem[112]=8'b0000000_0;
// mem[113]=8'b0101_0000;
// mem[114]=8'b0_010_0110;
// mem[115]=8'b0_0100011; //sw x5, 12(x0)
// mem[116]=8'b0000000_0;
// mem[117]=8'b0000_0000;
// mem[118]=8'b0_000_0000;
// mem[119]=8'b0_0110011 ; //add x0, x0, x0
// mem[120]=8'b0000000_0;
// mem[121]=8'b0000_0000;
// mem[122]=8'b0_000_0000;
// mem[123]=8'b0_0110011 ; //add x0, x0, x0
// mem[124]=8'b0000000_0;
// mem[125]=8'b0000_0000;
// mem[126]=8'b0_000_0000;
// mem[127]=8'b0_0110011 ; //add x0, x0, x0
// mem[128]=8'b00000000;
// mem[129]=8'b1100_0000;
// mem[130]=8'b0_010_0011;
// mem[131]=8'b0_0000011 ; //lw x6, 12(x0)
// mem[132]=8'b0000000_0;
// mem[133]=8'b0000_0000;
// mem[134]=8'b0_000_0000;
// mem[135]=8'b0_0110011 ; //add x0, x0, x0
// mem[136]=8'b0000000_0;
// mem[137]=8'b0000_0000;
// mem[138]=8'b0_000_0000;
// mem[139]=8'b0_0110011 ; //add x0, x0, x0
// mem[140]=8'b0000000_0;
// mem[141]=8'b0000_0000;
// mem[142]=8'b0_000_0000;
// mem[143]=8'b0_0110011 ; //add x0, x0, x0
// mem[144]=8'b0000000_0;
// mem[145]=8'b0001_0011;
// mem[146]=8'b0_111_0011;
// mem[147]=8'b1_0110011 ; //and x7, x6, x1
// mem[148]=8'b0000000_0;
// mem[149]=8'b0000_0000;
// mem[150]=8'b0_000_0000;
// mem[151]=8'b0_0110011 ; //add x0, x0, x0
// mem[152]=8'b0000000_0;
// mem[153]=8'b0000_0000;
// mem[154]=8'b0_000_0000;
// mem[155]=8'b0_0110011 ; //add x0, x0, x0
// mem[156]=8'b0000000_0;
// mem[157]=8'b0000_0000;
// mem[158]=8'b0_000_0000;
// mem[159]=8'b0_0110011 ; //add x0, x0, x0
// mem[160]=8'b0100000_0;
// mem[161]=8'b0010_0000;
// mem[162]=8'b1_000_0100;
// mem[163]=8'b0_0110011 ; //sub x8, x1, x2
// mem[164]=8'b0000000_0;
// mem[165]=8'b0000_0000;
// mem[166]=8'b0_000_0000;
// mem[167]=8'b0_0110011 ; //add x0, x0, x0
// mem[168]=8'b0000000_0;
// mem[169]=8'b0000_0000;
// mem[170]=8'b0_000_0000;
// mem[171]=8'b0_0110011 ; //add x0, x0, x0
// mem[172]=8'b0000000_0;
// mem[173]=8'b0000_0000;
// mem[174]=8'b0_000_0000;
// mem[175]=8'b0_0110011 ; //add x0, x0, x0
// mem[176]=8'b0000000_0;
// mem[177]=8'b0010_0000;
// mem[178]=8'b1_000_0000;
// mem[179]=8'b0_0110011 ; //add x0, x1, x2
// mem[180]=8'b0000000_0;
// mem[181]=8'b0000_0000;
// mem[182]=8'b0_000_0000;
// mem[183]=8'b0_0110011 ; //add x0, x0, x0
// mem[184]=8'b0000000_0;
// mem[185]=8'b0000_0000;
// mem[186]=8'b0_000_0000;
// mem[187]=8'b0_0110011 ; //add x0, x0, x0
// mem[188]=8'b0000000_0;
// mem[189]=8'b0000_0000;
// mem[190]=8'b0_000_0000;
// mem[191]=8'b0_0110011 ; //add x0, x0, x0
// mem[192]=8'b0000000_0;
// mem[193]=8'b0001_0000;
// mem[194]=8'b0_000_0100;
// mem[195]=8'b1_0110011 ; //add x9, x0, x1
//  end
//  mem[0]= 8'h00;
//  mem[1]= 8'h00;
//  mem[2]= 8'h24;
//  mem[3]= 8'h03;
  
//  mem[4]= 8'h00;
//  mem[5]= 8'h40;
//  mem[6]= 8'h24;
//  mem[7]= 8'h83;
  
//  mem[8]= 8'h00;
//  mem[9]= 8'h80;
//  mem[10]= 8'h21;
//  mem[11]= 8'h83;
  
//  mem[12]= 8'h00;
//  mem[13]= 8'h94;
//  mem[14]= 8'h65;
//  mem[15]= 8'h33;
  
//  mem[16]= 8'h00;
//  mem[17]= 8'h55;
//  mem[18]= 8'h05;
//  mem[19]= 8'h93;
  
//  mem[20]= 8'h00;
//  mem[21]= 8'h15;
//  mem[22]= 8'hd6;
//  mem[23]= 8'h13;
//  mem[24]= 8'h00;
//  mem[25]= 8'hc5;
//  mem[26]= 8'h21;
//  mem[27]= 8'h23;
//  mem[28]= 8'h00;
//  mem[29]= 8'h25;
//  mem[30]= 8'h27;
//  mem[31]= 8'h03;
//  mem[8]= 8'h00;
//  mem[33]= 8'hb7;
//  mem[34]= 8'h37;
//  mem[35]= 8'hb3;
  
// mem[36]= 8'hff;
// mem[37]= 8'hf7;
// mem[38]= 8'h26;
// mem[39]= 8'h93;
// mem[40]= 8'h25;
// mem[41]= 8'h80;
// mem[42]= 8'h00;
// mem[43]= 8'h93;
  
  
//  mem[44]= 8'h00;
//  mem[45]= 8'h15;
//  mem[46]= 8'h20;
//  mem[47]= 8'h23;
  
//  mem[48]= 8'h00;
//    mem[49]= 8'h05;
//    mem[50]= 8'h08;
//    mem[51]= 8'h03;
//    mem[52]= 8'h00;
//      mem[53]= 8'h85;
//      mem[54]= 8'h11;
//      mem[55]= 8'h33;
//      mem[56]= 8'h00;
//        mem[57]= 8'h10;
//        mem[58]= 8'h00;
//        mem[59]= 8'h73;
  
//  end 

 
 
 
//initial begin


//end
 assign instruction = {mem[address],mem[address+1],mem[address+2],mem[((address)+3)]}; 
     
endmodule
